module testbench();
    reg clk;
    reg rst;
    
    soc_top u_soc_top(
    	.clk (clk ),
        .rst (rst )
    );
    

    initial begin
        clk = 1'b0;
        rst = 1'b0;
        // rom[0] = 31'b00111100000000010000000000000001;
        // rom[1] = 31'b00000000000000010000100001000000;
        // rom[2] = 31'b00010000000000000000000000000100;
        // rom[3] = 31'b00000000000000010000100001000000;
        // rom[4] = 31'b00000000000000010000100001000000;
        // rom[5] = 31'b00000000000000010000100001000000;
        // rom[6] = 31'b00000000000000010000100001000000;
        // rom[7] = 31'b00000000000000010000100001000000;
        #10
        rst = 1'b1;
        #30
        rst = 1'b0;    
    end

    always # 5 clk = ~clk;
    // always @ (*) begin
    //     inst = rom[inst_addr[4:2]];
    // end

endmodule 