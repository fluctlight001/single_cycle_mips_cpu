`include "defines.vh"
module rom(
    input wire clk,
    input wire rst,
    input wire [31:0] addr,
    output reg [31:0] data
);
    reg [31:0] rom [7:0];
    always @ (posedge clk) begin
        if (rst == `RstEnable) begin
            // rom[0] <= 31'b00111100000000010000000000000001;
            // rom[1] <= 31'b00000000000000010000100001000000;
            // rom[2] <= 31'b00010000000000000000000000000100;
            // rom[3] <= 31'b00000000000000010000100001000000;
            // rom[4] <= 31'b00000000000000010000100001000000;
            // rom[5] <= 31'b00000000000000010000100001000000;
            // rom[6] <= 31'b00000000000000010000100001000000;
            // rom[7] <= 31'b00000000000000010000100001000000;
            rom[0] <= 32'b00111100000000010000000000000001;
            rom[1] <= 32'b00111100000000100000000000000001;
            rom[2] <= 32'b00000000001000100000100000100001;
            rom[3] <= 32'b00000000001000100001000000100001;
            rom[4] <= 32'b10101100000000100000000000000000;
            rom[5] <= 32'b10001100000000110000000000000000;
            rom[6] <= 32'b00111100000001000000000000000011;
            rom[7] <= 32'b00010000011001000000000000001000;
            // command
            // LUI 1 1
            // LUI 2 1
            // ADDU 1 1 2
            // ADDU 2 1 2
            // SW 2 0 0
            // LW 3 0 0
            // LUI 4 3
            // BEQ 3 4 8
        end
    end
    always @ (*) begin
        data = rom[addr[4:2]];
    end
endmodule 